`timescale 1ns / 1ps
//*************************************************************************
//   > �ļ���: single_cycle_cpu.v
//   > ����  :������CPUģ�飬��ʵ��16��ָ��
//   >        ָ��rom������ram�������첽�����ݣ��Ա㵥����CPU��ʵ��
//   > ����  : LOONGSON
//   > ����  : 2016-04-14
//*************************************************************************
`define STARTADDR 32'd0 
module single_cycle_cpu(
    input clk,   
    input resetn, 

    input  [ 4:0] rf_addr,
    input  [31:0] mem_addr,
    output [31:0] rf_data,
    output [31:0] mem_data,
    output [31:0] cpu_pc,
    output [31:0] cpu_inst
    );

//---------------------------------{ȡָ}begin------------------------------------//

//���ڴ˴���Ӵ���

//----------------------------------{ȡָ}end-------------------------------------//

//---------------------------------{����}begin------------------------------------//

//���ڴ˴���Ӵ���

//----------------------------------{����}end-------------------------------------//

//---------------------------------{ִ��}begin------------------------------------//

//���ڴ˴���Ӵ���

//----------------------------------{ִ��}end-------------------------------------//
    
//---------------------------------{�ô�}begin------------------------------------//

//���ڴ˴���Ӵ���

//----------------------------------{�ô�}end-------------------------------------//

//---------------------------------{д��}begin------------------------------------//

//���ڴ˴���Ӵ���

//----------------------------------{д��}end-------------------------------------//
endmodule
